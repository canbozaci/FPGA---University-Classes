`timescale 1ns / 1ps

module SSI_Library(

    );

endmodule 
// ----------  ----------  ----------  ----------  	OR_GATE	   ----------  ----------  ----------  ---------- 
module OR(
	output O,
	input I1,
	input I2
    );
	assign O = I1 | I2;
endmodule
// ----------  ----------  ----------  ----------  ----------  ----------  ----------  ----------  ---------- 

// ----------  ----------  ----------  ----------  	NOT_GATE   ----------  ----------  ----------  ---------- 
module NOT(
	output O,
	input I
    );
	assign O = ~I;
endmodule
// ----------  ----------  ----------  ----------  ----------  ----------  ----------  ----------  ---------- 


// ----------  ----------  ----------  ----------  	NAND_GATE  ----------  ----------  ----------  ---------- 
module NAND(
	output reg O,
	input I1,
	input I2
    );
	always@(*)
	begin
	O=~(I1 & I2);
	end
endmodule
// ----------  ----------  ----------  ----------  ----------  ----------  ----------  ----------  ---------- 

// ----------  ----------  ----------  ----------  	NOR_GATE   ----------  ----------  ----------  ---------- 
module NOR(
	output reg O,
	input I1,
	input I2
    );
	always@(*)
	begin
	O=~(I1 | I2);
	end
endmodule
// ----------  ----------  ----------  ----------  ----------  ----------  ----------  ----------  ---------- 

// ----------  ----------  ----------  ----------  	EXOR_GATE  ----------  ----------  ----------  ---------- 
module EXOR(
	output O,
	input I1,
	input I2
    );
	LUT2#(.INIT(4'b0110))lut(.O(O),.I1(I1),.I0(I2));
endmodule
// ----------  ----------  ----------  ----------  ----------  ----------  ----------  ----------  ----------

// ----------  ----------  ----------  ----------  	EXNOR_GATE ----------  ----------  ----------  ---------- 
module EXNOR(
	output O,
	input I1,
	input I2
    );
	LUT2#(.INIT(4'b1001))lut(.O(O),.I1(I1),.I0(I2));
endmodule
// ----------  ----------  ----------  ----------  ----------  ----------  ----------  ----------  ---------- 

// ----------  ----------  ----------  ----------  TRI_GATE	   ----------  ----------  ----------  ---------- 
module TRI(
	output O,
	input I,
	input E
    );
	assign O = E ? I : 1'bz;
endmodule
// ----------  ----------  ----------  ----------  ----------  ----------  ----------  ----------  ---------- 

// ----------  ----------  ----------  ----------  TOP_MODULE  ----------  ----------  ----------  ---------- 
/*module TOP(
output O_or,
output O_not,
output O_nand,
output O_nor,
output O_exor,
output O_exnor,
output O_tri,
input I1,
input I2
    );

OR or_gate(O_or, I1, I2);
NOT not_gate(O_not, I1);
NAND nand_gate(O_nand,I1,I2);
NOR nor_gate(O_nor,I1,I2);
EXOR exor_gate(O_exor,I1,I2);
EXNOR exnor_gate(O_exnor,I1,I2);
TRI tri_gate(O_tri,I1,I2);


endmodule*/
// ----------  ----------  ----------  ----------  ----------  ----------  ----------  ----------  ---------- 