`timescale 1ns / 1ps
module arccosh(
	input [10:0] x,
	output reg [7:0] y
    );
always@(*) begin
	case(x)
	11'b00000100000  : y = 8'b00000000 ;
    11'b00000100001  : y = 8'b00000011 ;
	11'b00000100010  : y = 8'b00000101 ;
    11'b00000100011  : y = 8'b00000110 ;
	11'b00000100100  : y = 8'b00000111 ;
	11'b00000100101  : y = 8'b00001000 ;
	11'b00000100110  : y = 8'b00001001 ;
	11'b00000100111  : y = 8'b00001010 ;
	11'b00000101000  : y = 8'b00001011 ;
    11'b00000101001  : y = 8'b00001011 ;
    11'b00000101010  : y = 8'b00001100 ;
    11'b00000101011  : y = 8'b00001100 ;
    11'b00000101100  : y = 8'b00001101 ;
    11'b00000101101  : y = 8'b00001101 ;
    11'b00000101110  : y = 8'b00001110 ;
    11'b00000101111  : y = 8'b00001110 ;
    11'b00000110000  : y = 8'b00001111 ;
    11'b00000110001  : y = 8'b00001111 ;
    11'b00000110010  : y = 8'b00010000 ;
    11'b00000110011  : y = 8'b00010000 ;
    11'b00000110100  : y = 8'b00010001 ;
    11'b00000110101  : y = 8'b00010001 ;
    11'b00000110110  : y = 8'b00010001 ;
    11'b00000110111  : y = 8'b00010010 ;
    11'b00000111000  : y = 8'b00010010 ;
    11'b00000111001  : y = 8'b00010010 ;
    11'b00000111010  : y = 8'b00010011 ;
    11'b00000111011  : y = 8'b00010011 ;
    11'b00000111100  : y = 8'b00010011 ;
    11'b00000111101  : y = 8'b00010100 ;
    11'b00000111110  : y = 8'b00010100 ;
    11'b00000111111  : y = 8'b00010100 ;
    11'b00001000000  : y = 8'b00010101 ;
    11'b00001000001  : y = 8'b00010101 ;
    11'b00001000010  : y = 8'b00010101 ;
    11'b00001000011  : y = 8'b00010101 ;
    11'b00001000100  : y = 8'b00010110 ;
    11'b00001000101  : y = 8'b00010110 ;
    11'b00001000110  : y = 8'b00010110 ;
    11'b00001000111  : y = 8'b00010110 ;
    11'b00001001000  : y = 8'b00010111 ;
    11'b00001001001  : y = 8'b00010111 ;
    11'b00001001010  : y = 8'b00010111 ;
    11'b00001001011  : y = 8'b00010111 ;
    11'b00001001100  : y = 8'b00011000 ;
    11'b00001001101  : y = 8'b00011000 ;
    11'b00001001110  : y = 8'b00011000 ;
    11'b00001001111  : y = 8'b00011000 ;
    11'b00001010000  : y = 8'b00011001 ;
    11'b00001010001  : y = 8'b00011001 ;
    11'b00001010010  : y = 8'b00011001 ;
    11'b00001010011  : y = 8'b00011001 ;
    11'b00001010100  : y = 8'b00011001 ;
    11'b00001010101  : y = 8'b00011010 ;
    11'b00001010110  : y = 8'b00011010 ;
    11'b00001010111  : y = 8'b00011010 ;
    11'b00001011000  : y = 8'b00011010 ;
    11'b00001011001  : y = 8'b00011010 ;
    11'b00001011010  : y = 8'b00011011 ;
    11'b00001011011  : y = 8'b00011011 ;
    11'b00001011100  : y = 8'b00011011 ;
    11'b00001011101  : y = 8'b00011011 ;
    11'b00001011110  : y = 8'b00011011 ;
    11'b00001011111  : y = 8'b00011100 ;
    11'b00001100000  : y = 8'b00011100 ;
    11'b00001100001  : y = 8'b00011100 ;
    11'b00001100010  : y = 8'b00011100 ;
    11'b00001100011  : y = 8'b00011100 ;
    11'b00001100100  : y = 8'b00011100 ;
    11'b00001100101  : y = 8'b00011101 ;
    11'b00001100110  : y = 8'b00011101 ;
    11'b00001100111  : y = 8'b00011101 ;
    11'b00001101000  : y = 8'b00011101 ;
    11'b00001101001  : y = 8'b00011101 ;
    11'b00001101010  : y = 8'b00011101 ;
    11'b00001101011  : y = 8'b00011110 ;
    11'b00001101100  : y = 8'b00011110 ;
    11'b00001101101  : y = 8'b00011110 ;
    11'b00001101110  : y = 8'b00011110 ;
    11'b00001101111  : y = 8'b00011110 ;
    11'b00001110000  : y = 8'b00011110 ;
    11'b00001110001  : y = 8'b00011110 ;
    11'b00001110010  : y = 8'b00011111 ;
    11'b00001110011  : y = 8'b00011111 ;
    11'b00001110100  : y = 8'b00011111 ;
    11'b00001110101  : y = 8'b00011111 ;
    11'b00001110110  : y = 8'b00011111 ;
    11'b00001110111  : y = 8'b00011111 ;
    11'b00001111000  : y = 8'b00011111 ;
    11'b00001111001  : y = 8'b00100000 ;
    11'b00001111010  : y = 8'b00100000 ;
    11'b00001111011  : y = 8'b00100000 ;
    11'b00001111100  : y = 8'b00100000 ;
    11'b00001111101  : y = 8'b00100000 ;
    11'b00001111110  : y = 8'b00100000 ;
    11'b00001111111  : y = 8'b00100000 ;
    11'b00010000000  : y = 8'b00100001 ;
    11'b00010000001  : y = 8'b00100001 ;
    11'b00010000010  : y = 8'b00100001 ;
    11'b00010000011  : y = 8'b00100001 ;
    11'b00010000100  : y = 8'b00100001 ;
    11'b00010000101  : y = 8'b00100001 ;
    11'b00010000110  : y = 8'b00100001 ;
    11'b00010000111  : y = 8'b00100001 ;
    11'b00010001000  : y = 8'b00100010 ;
    11'b00010001001  : y = 8'b00100010 ;
    11'b00010001010  : y = 8'b00100010 ;
    11'b00010001011  : y = 8'b00100010 ;
    11'b00010001100  : y = 8'b00100010 ;
    11'b00010001101  : y = 8'b00100010 ;
    11'b00010001110  : y = 8'b00100010 ;
    11'b00010001111  : y = 8'b00100010 ;
    11'b00010010000  : y = 8'b00100010 ;
    11'b00010010001  : y = 8'b00100011 ;
    11'b00010010010  : y = 8'b00100011 ;
    11'b00010010011  : y = 8'b00100011 ;
    11'b00010010100  : y = 8'b00100011 ;
    11'b00010010101  : y = 8'b00100011 ;
    11'b00010010110  : y = 8'b00100011 ;
    11'b00010010111  : y = 8'b00100011 ;
    11'b00010011000  : y = 8'b00100011 ;
    11'b00010011001  : y = 8'b00100011 ;
    11'b00010011010  : y = 8'b00100100 ;
    11'b00010011011  : y = 8'b00100100 ;
    11'b00010011100  : y = 8'b00100100 ;
    11'b00010011101  : y = 8'b00100100 ;
    11'b00010011110  : y = 8'b00100100 ;
    11'b00010011111  : y = 8'b00100100 ;
    11'b00010100000  : y = 8'b00100100 ;
    11'b00010100001  : y = 8'b00100100 ;
    11'b00010100010  : y = 8'b00100100 ;
    11'b00010100011  : y = 8'b00100100 ;
    11'b00010100100  : y = 8'b00100101 ;
    11'b00010100101  : y = 8'b00100101 ;
    11'b00010100110  : y = 8'b00100101 ;
    11'b00010100111  : y = 8'b00100101 ;
    11'b00010101000  : y = 8'b00100101 ;
    11'b00010101001  : y = 8'b00100101 ;
    11'b00010101010  : y = 8'b00100101 ;
    11'b00010101011  : y = 8'b00100101 ;
    11'b00010101100  : y = 8'b00100101 ;
    11'b00010101101  : y = 8'b00100101 ;
    11'b00010101110  : y = 8'b00100110 ;
    11'b00010101111  : y = 8'b00100110 ;
    11'b00010110000  : y = 8'b00100110 ;
    11'b00010110001  : y = 8'b00100110 ;
    11'b00010110010  : y = 8'b00100110 ;
    11'b00010110011  : y = 8'b00100110 ;
    11'b00010110100  : y = 8'b00100110 ;
    11'b00010110101  : y = 8'b00100110 ;
    11'b00010110110  : y = 8'b00100110 ;
    11'b00010110111  : y = 8'b00100110 ;
    11'b00010111000  : y = 8'b00100110 ;
    11'b00010111001  : y = 8'b00100111 ;
    11'b00010111010  : y = 8'b00100111 ;
    11'b00010111011  : y = 8'b00100111 ;
    11'b00010111100  : y = 8'b00100111 ;
    11'b00010111101  : y = 8'b00100111 ;
    11'b00010111110  : y = 8'b00100111 ;
    11'b00010111111  : y = 8'b00100111 ;
    11'b00011000000  : y = 8'b00100111 ;
    11'b00011000001  : y = 8'b00100111 ;
    11'b00011000010  : y = 8'b00100111 ;
    11'b00011000011  : y = 8'b00100111 ;
    11'b00011000100  : y = 8'b00100111 ;
    11'b00011000101  : y = 8'b00101000 ;
    11'b00011000110  : y = 8'b00101000 ;
    11'b00011000111  : y = 8'b00101000 ;
    11'b00011001000  : y = 8'b00101000 ;
    11'b00011001001  : y = 8'b00101000 ;
    11'b00011001010  : y = 8'b00101000 ;
    11'b00011001011  : y = 8'b00101000 ;
    11'b00011001100  : y = 8'b00101000 ;
    11'b00011001101  : y = 8'b00101000 ;
    11'b00011001110  : y = 8'b00101000 ;
    11'b00011001111  : y = 8'b00101000 ;
    11'b00011010000  : y = 8'b00101000 ;
    11'b00011010001  : y = 8'b00101001 ;
    11'b00011010010  : y = 8'b00101001 ;
    11'b00011010011  : y = 8'b00101001 ;
    11'b00011010100  : y = 8'b00101001 ;
    11'b00011010101  : y = 8'b00101001 ;
    11'b00011010110  : y = 8'b00101001 ;
    11'b00011010111  : y = 8'b00101001 ;
    11'b00011011000  : y = 8'b00101001 ;
    11'b00011011001  : y = 8'b00101001 ;
    11'b00011011010  : y = 8'b00101001 ;
    11'b00011011011  : y = 8'b00101001 ;
    11'b00011011100  : y = 8'b00101001 ;
    11'b00011011101  : y = 8'b00101001 ;
    11'b00011011110  : y = 8'b00101001 ;
    11'b00011011111  : y = 8'b00101010 ;
    11'b00011100000  : y = 8'b00101010 ;
    11'b00011100001  : y = 8'b00101010 ;
    11'b00011100010  : y = 8'b00101010 ;
    11'b00011100011  : y = 8'b00101010 ;
    11'b00011100100  : y = 8'b00101010 ;
    11'b00011100101  : y = 8'b00101010 ;
    11'b00011100110  : y = 8'b00101010 ;
    11'b00011100111  : y = 8'b00101010 ;
    11'b00011101000  : y = 8'b00101010 ;
    11'b00011101001  : y = 8'b00101010 ;
    11'b00011101010  : y = 8'b00101010 ;
    11'b00011101011  : y = 8'b00101010 ;
    11'b00011101100  : y = 8'b00101010 ;
    11'b00011101101  : y = 8'b00101011 ;
    11'b00011101110  : y = 8'b00101011 ;
    11'b00011101111  : y = 8'b00101011 ;
    11'b00011110000  : y = 8'b00101011 ;
    11'b00011110001  : y = 8'b00101011 ;
    11'b00011110010  : y = 8'b00101011 ;
    11'b00011110011  : y = 8'b00101011 ;
    11'b00011110100  : y = 8'b00101011 ;
    11'b00011110101  : y = 8'b00101011 ;
    11'b00011110110  : y = 8'b00101011 ;
    11'b00011110111  : y = 8'b00101011 ;
    11'b00011111000  : y = 8'b00101011 ;
    11'b00011111001  : y = 8'b00101011 ;
    11'b00011111010  : y = 8'b00101011 ;
    11'b00011111011  : y = 8'b00101011 ;
    11'b00011111100  : y = 8'b00101100 ;
    11'b00011111101  : y = 8'b00101100 ;
    11'b00011111110  : y = 8'b00101100 ;
    11'b00011111111  : y = 8'b00101100 ;
    11'b00100000000  : y = 8'b00101100 ;
    11'b00100000001  : y = 8'b00101100 ;
    11'b00100000010  : y = 8'b00101100 ;
    11'b00100000011  : y = 8'b00101100 ;
    11'b00100000100  : y = 8'b00101100 ;
    11'b00100000101  : y = 8'b00101100 ;
    11'b00100000110  : y = 8'b00101100 ;
    11'b00100000111  : y = 8'b00101100 ;
    11'b00100001000  : y = 8'b00101100 ;
    11'b00100001001  : y = 8'b00101100 ;
    11'b00100001010  : y = 8'b00101100 ;
    11'b00100001011  : y = 8'b00101100 ;
    11'b00100001100  : y = 8'b00101101 ;
    11'b00100001101  : y = 8'b00101101 ;
    11'b00100001110  : y = 8'b00101101 ;
    11'b00100001111  : y = 8'b00101101 ;
    11'b00100010000  : y = 8'b00101101 ;
    11'b00100010001  : y = 8'b00101101 ;
    11'b00100010010  : y = 8'b00101101 ;
    11'b00100010011  : y = 8'b00101101 ;
    11'b00100010100  : y = 8'b00101101 ;
    11'b00100010101  : y = 8'b00101101 ;
    11'b00100010110  : y = 8'b00101101 ;
    11'b00100010111  : y = 8'b00101101 ;
    11'b00100011000  : y = 8'b00101101 ;
    11'b00100011001  : y = 8'b00101101 ;
    11'b00100011010  : y = 8'b00101101 ;
    11'b00100011011  : y = 8'b00101101 ;
    11'b00100011100  : y = 8'b00101101 ;
    11'b00100011101  : y = 8'b00101110 ;
    11'b00100011110  : y = 8'b00101110 ;
    11'b00100011111  : y = 8'b00101110 ;
    11'b00100100000  : y = 8'b00101110 ;
    11'b00100100001  : y = 8'b00101110 ;
    11'b00100100010  : y = 8'b00101110 ;
    11'b00100100011  : y = 8'b00101110 ;
    11'b00100100100  : y = 8'b00101110 ;
    11'b00100100101  : y = 8'b00101110 ;
    11'b00100100110  : y = 8'b00101110 ;
    11'b00100100111  : y = 8'b00101110 ;
    11'b00100101000  : y = 8'b00101110 ;
    11'b00100101001  : y = 8'b00101110 ;
    11'b00100101010  : y = 8'b00101110 ;
    11'b00100101011  : y = 8'b00101110 ;
    11'b00100101100  : y = 8'b00101110 ;
    11'b00100101101  : y = 8'b00101110 ;
    11'b00100101110  : y = 8'b00101110 ;
    11'b00100101111  : y = 8'b00101111 ;
    11'b00100110000  : y = 8'b00101111 ;
    11'b00100110001  : y = 8'b00101111 ;
    11'b00100110010  : y = 8'b00101111 ;
    11'b00100110011  : y = 8'b00101111 ;
    11'b00100110100  : y = 8'b00101111 ;
    11'b00100110101  : y = 8'b00101111 ;
    11'b00100110110  : y = 8'b00101111 ;
    11'b00100110111  : y = 8'b00101111 ;
    11'b00100111000  : y = 8'b00101111 ;
    11'b00100111001  : y = 8'b00101111 ;
    11'b00100111010  : y = 8'b00101111 ;
    11'b00100111011  : y = 8'b00101111 ;
    11'b00100111100  : y = 8'b00101111 ;
    11'b00100111101  : y = 8'b00101111 ;
    11'b00100111110  : y = 8'b00101111 ;
    11'b00100111111  : y = 8'b00101111 ;
    11'b00101000000  : y = 8'b00101111 ;
    11'b00101000001  : y = 8'b00101111 ;
    11'b00101000010  : y = 8'b00101111 ;
    11'b00101000011  : y = 8'b00110000 ;
    11'b00101000100  : y = 8'b00110000 ;
    11'b00101000101  : y = 8'b00110000 ;
    11'b00101000110  : y = 8'b00110000 ;
    11'b00101000111  : y = 8'b00110000 ;
    11'b00101001000  : y = 8'b00110000 ;
    11'b00101001001  : y = 8'b00110000 ;
    11'b00101001010  : y = 8'b00110000 ;
    11'b00101001011  : y = 8'b00110000 ;
    11'b00101001100  : y = 8'b00110000 ;
    11'b00101001101  : y = 8'b00110000 ;
    11'b00101001110  : y = 8'b00110000 ;
    11'b00101001111  : y = 8'b00110000 ;
    11'b00101010000  : y = 8'b00110000 ;
    11'b00101010001  : y = 8'b00110000 ;
    11'b00101010010  : y = 8'b00110000 ;
    11'b00101010011  : y = 8'b00110000 ;
    11'b00101010100  : y = 8'b00110000 ;
    11'b00101010101  : y = 8'b00110000 ;
    11'b00101010110  : y = 8'b00110000 ;
    11'b00101010111  : y = 8'b00110001 ;
    11'b00101011000  : y = 8'b00110001 ;
    11'b00101011001  : y = 8'b00110001 ;
    11'b00101011010  : y = 8'b00110001 ;
    11'b00101011011  : y = 8'b00110001 ;
    11'b00101011100  : y = 8'b00110001 ;
    11'b00101011101  : y = 8'b00110001 ;
    11'b00101011110  : y = 8'b00110001 ;
    11'b00101011111  : y = 8'b00110001 ;
    11'b00101100000  : y = 8'b00110001 ;
    11'b00101100001  : y = 8'b00110001 ;
    11'b00101100010  : y = 8'b00110001 ;
    11'b00101100011  : y = 8'b00110001 ;
    11'b00101100100  : y = 8'b00110001 ;
    11'b00101100101  : y = 8'b00110001 ;
    11'b00101100110  : y = 8'b00110001 ;
    11'b00101100111  : y = 8'b00110001 ;
    11'b00101101000  : y = 8'b00110001 ;
    11'b00101101001  : y = 8'b00110001 ;
    11'b00101101010  : y = 8'b00110001 ;
    11'b00101101011  : y = 8'b00110001 ;
    11'b00101101100  : y = 8'b00110001 ;
    11'b00101101101  : y = 8'b00110010 ;
    11'b00101101110  : y = 8'b00110010 ;
    11'b00101101111  : y = 8'b00110010 ;
    11'b00101110000  : y = 8'b00110010 ;
    11'b00101110001  : y = 8'b00110010 ;
    11'b00101110010  : y = 8'b00110010 ;
    11'b00101110011  : y = 8'b00110010 ;
    11'b00101110100  : y = 8'b00110010 ;
    11'b00101110101  : y = 8'b00110010 ;
    11'b00101110110  : y = 8'b00110010 ;
    11'b00101110111  : y = 8'b00110010 ;
    11'b00101111000  : y = 8'b00110010 ;
    11'b00101111001  : y = 8'b00110010 ;
    11'b00101111010  : y = 8'b00110010 ;
    11'b00101111011  : y = 8'b00110010 ;
    11'b00101111100  : y = 8'b00110010 ;
    11'b00101111101  : y = 8'b00110010 ;
    11'b00101111110  : y = 8'b00110010 ;
    11'b00101111111  : y = 8'b00110010 ;
    11'b00110000000  : y = 8'b00110010 ;
    11'b00110000001  : y = 8'b00110010 ;
    11'b00110000010  : y = 8'b00110010 ;
    11'b00110000011  : y = 8'b00110010 ;
    11'b00110000100  : y = 8'b00110010 ;
    11'b00110000101  : y = 8'b00110011 ;
    11'b00110000110  : y = 8'b00110011 ;
    11'b00110000111  : y = 8'b00110011 ;
    11'b00110001000  : y = 8'b00110011 ;
    11'b00110001001  : y = 8'b00110011 ;
    11'b00110001010  : y = 8'b00110011 ;
    11'b00110001011  : y = 8'b00110011 ;
    11'b00110001100  : y = 8'b00110011 ;
    11'b00110001101  : y = 8'b00110011 ;
    11'b00110001110  : y = 8'b00110011 ;
    11'b00110001111  : y = 8'b00110011 ;
    11'b00110010000  : y = 8'b00110011 ;
    11'b00110010001  : y = 8'b00110011 ;
    11'b00110010010  : y = 8'b00110011 ;
    11'b00110010011  : y = 8'b00110011 ;
    11'b00110010100  : y = 8'b00110011 ;
    11'b00110010101  : y = 8'b00110011 ;
    11'b00110010110  : y = 8'b00110011 ;
    11'b00110010111  : y = 8'b00110011 ;
    11'b00110011000  : y = 8'b00110011 ;
    11'b00110011001  : y = 8'b00110011 ;
    11'b00110011010  : y = 8'b00110011 ;
    11'b00110011011  : y = 8'b00110011 ;
    11'b00110011100  : y = 8'b00110011 ;
    11'b00110011101  : y = 8'b00110011 ;
    11'b00110011110  : y = 8'b00110100 ;
    11'b00110011111  : y = 8'b00110100 ;
    11'b00110100000  : y = 8'b00110100 ;
    11'b00110100001  : y = 8'b00110100 ;
    11'b00110100010  : y = 8'b00110100 ;
    11'b00110100011  : y = 8'b00110100 ;
    11'b00110100100  : y = 8'b00110100 ;
    11'b00110100101  : y = 8'b00110100 ;
    11'b00110100110  : y = 8'b00110100 ;
    11'b00110100111  : y = 8'b00110100 ;
    11'b00110101000  : y = 8'b00110100 ;
    11'b00110101001  : y = 8'b00110100 ;
    11'b00110101010  : y = 8'b00110100 ;
    11'b00110101011  : y = 8'b00110100 ;
    11'b00110101100  : y = 8'b00110100 ;
    11'b00110101101  : y = 8'b00110100 ;
    11'b00110101110  : y = 8'b00110100 ;
    11'b00110101111  : y = 8'b00110100 ;
    11'b00110110000  : y = 8'b00110100 ;
    11'b00110110001  : y = 8'b00110100 ;
    11'b00110110010  : y = 8'b00110100 ;
    11'b00110110011  : y = 8'b00110100 ;
    11'b00110110100  : y = 8'b00110100 ;
    11'b00110110101  : y = 8'b00110100 ;
    11'b00110110110  : y = 8'b00110100 ;
    11'b00110110111  : y = 8'b00110100 ;
    11'b00110111000  : y = 8'b00110101 ;
    11'b00110111001  : y = 8'b00110101 ;
    11'b00110111010  : y = 8'b00110101 ;
    11'b00110111011  : y = 8'b00110101 ;
    11'b00110111100  : y = 8'b00110101 ;
    11'b00110111101  : y = 8'b00110101 ;
    11'b00110111110  : y = 8'b00110101 ;
    11'b00110111111  : y = 8'b00110101 ;
    11'b00111000000  : y = 8'b00110101 ;
    11'b00111000001  : y = 8'b00110101 ;
    11'b00111000010  : y = 8'b00110101 ;
    11'b00111000011  : y = 8'b00110101 ;
    11'b00111000100  : y = 8'b00110101 ;
    11'b00111000101  : y = 8'b00110101 ;
    11'b00111000110  : y = 8'b00110101 ;
    11'b00111000111  : y = 8'b00110101 ;
    11'b00111001000  : y = 8'b00110101 ;
    11'b00111001001  : y = 8'b00110101 ;
    11'b00111001010  : y = 8'b00110101 ;
    11'b00111001011  : y = 8'b00110101 ;
    11'b00111001100  : y = 8'b00110101 ;
    11'b00111001101  : y = 8'b00110101 ;
    11'b00111001110  : y = 8'b00110101 ;
    11'b00111001111  : y = 8'b00110101 ;
    11'b00111010000  : y = 8'b00110101 ;
    11'b00111010001  : y = 8'b00110101 ;
    11'b00111010010  : y = 8'b00110101 ;
    11'b00111010011  : y = 8'b00110101 ;
    11'b00111010100  : y = 8'b00110101 ;
    11'b00111010101  : y = 8'b00110110 ;
    11'b00111010110  : y = 8'b00110110 ;
    11'b00111010111  : y = 8'b00110110 ;
    11'b00111011000  : y = 8'b00110110 ;
    11'b00111011001  : y = 8'b00110110 ;
    11'b00111011010  : y = 8'b00110110 ;
    11'b00111011011  : y = 8'b00110110 ;
    11'b00111011100  : y = 8'b00110110 ;
    11'b00111011101  : y = 8'b00110110 ;
    11'b00111011110  : y = 8'b00110110 ;
    11'b00111011111  : y = 8'b00110110 ;
    11'b00111100000  : y = 8'b00110110 ;
    11'b00111100001  : y = 8'b00110110 ;
    11'b00111100010  : y = 8'b00110110 ;
    11'b00111100011  : y = 8'b00110110 ;
    11'b00111100100  : y = 8'b00110110 ;
    11'b00111100101  : y = 8'b00110110 ;
    11'b00111100110  : y = 8'b00110110 ;
    11'b00111100111  : y = 8'b00110110 ;
    11'b00111101000  : y = 8'b00110110 ;
    11'b00111101001  : y = 8'b00110110 ;
    11'b00111101010  : y = 8'b00110110 ;
    11'b00111101011  : y = 8'b00110110 ;
    11'b00111101100  : y = 8'b00110110 ;
    11'b00111101101  : y = 8'b00110110 ;
    11'b00111101110  : y = 8'b00110110 ;
    11'b00111101111  : y = 8'b00110110 ;
    11'b00111110000  : y = 8'b00110110 ;
    11'b00111110001  : y = 8'b00110110 ;
    11'b00111110010  : y = 8'b00110110 ;
    11'b00111110011  : y = 8'b00110111 ;
    11'b00111110100  : y = 8'b00110111 ;
    11'b00111110101  : y = 8'b00110111 ;
    11'b00111110110  : y = 8'b00110111 ;
    11'b00111110111  : y = 8'b00110111 ;
    11'b00111111000  : y = 8'b00110111 ;
    11'b00111111001  : y = 8'b00110111 ;
    11'b00111111010  : y = 8'b00110111 ;
    11'b00111111011  : y = 8'b00110111 ;
    11'b00111111100  : y = 8'b00110111 ;
    11'b00111111101  : y = 8'b00110111 ;
    11'b00111111110  : y = 8'b00110111 ;
    11'b00111111111  : y = 8'b00110111 ;
    11'b01000000000  : y = 8'b00110111 ;
    11'b01000000001  : y = 8'b00110111 ;
    11'b01000000010  : y = 8'b00110111 ;
    11'b01000000011  : y = 8'b00110111 ;
    11'b01000000100  : y = 8'b00110111 ;
    11'b01000000101  : y = 8'b00110111 ;
    11'b01000000110  : y = 8'b00110111 ;
    11'b01000000111  : y = 8'b00110111 ;
    11'b01000001000  : y = 8'b00110111 ;
    11'b01000001001  : y = 8'b00110111 ;
    11'b01000001010  : y = 8'b00110111 ;
    11'b01000001011  : y = 8'b00110111 ;
    11'b01000001100  : y = 8'b00110111 ;
    11'b01000001101  : y = 8'b00110111 ;
    11'b01000001110  : y = 8'b00110111 ;
    11'b01000001111  : y = 8'b00110111 ;
    11'b01000010000  : y = 8'b00110111 ;
    11'b01000010001  : y = 8'b00110111 ;
    11'b01000010010  : y = 8'b00110111 ;
    11'b01000010011  : y = 8'b00111000 ;
    11'b01000010100  : y = 8'b00111000 ;
    11'b01000010101  : y = 8'b00111000 ;
    11'b01000010110  : y = 8'b00111000 ;
    11'b01000010111  : y = 8'b00111000 ;
    11'b01000011000  : y = 8'b00111000 ;
    11'b01000011001  : y = 8'b00111000 ;
    11'b01000011010  : y = 8'b00111000 ;
    11'b01000011011  : y = 8'b00111000 ;
    11'b01000011100  : y = 8'b00111000 ;
    11'b01000011101  : y = 8'b00111000 ;
    11'b01000011110  : y = 8'b00111000 ;
    11'b01000011111  : y = 8'b00111000 ;
    11'b01000100000  : y = 8'b00111000 ;
    11'b01000100001  : y = 8'b00111000 ;
    11'b01000100010  : y = 8'b00111000 ;
    11'b01000100011  : y = 8'b00111000 ;
    11'b01000100100  : y = 8'b00111000 ;
    11'b01000100101  : y = 8'b00111000 ;
    11'b01000100110  : y = 8'b00111000 ;
    11'b01000100111  : y = 8'b00111000 ;
    11'b01000101000  : y = 8'b00111000 ;
    11'b01000101001  : y = 8'b00111000 ;
    11'b01000101010  : y = 8'b00111000 ;
    11'b01000101011  : y = 8'b00111000 ;
    11'b01000101100  : y = 8'b00111000 ;
    11'b01000101101  : y = 8'b00111000 ;
    11'b01000101110  : y = 8'b00111000 ;
    11'b01000101111  : y = 8'b00111000 ;
    11'b01000110000  : y = 8'b00111000 ;
    11'b01000110001  : y = 8'b00111000 ;
    11'b01000110010  : y = 8'b00111000 ;
    11'b01000110011  : y = 8'b00111000 ;
    11'b01000110100  : y = 8'b00111000 ;
    11'b01000110101  : y = 8'b00111001 ;
    11'b01000110110  : y = 8'b00111001 ;
    11'b01000110111  : y = 8'b00111001 ;
    11'b01000111000  : y = 8'b00111001 ;
    11'b01000111001  : y = 8'b00111001 ;
    11'b01000111010  : y = 8'b00111001 ;
    11'b01000111011  : y = 8'b00111001 ;
    11'b01000111100  : y = 8'b00111001 ;
    11'b01000111101  : y = 8'b00111001 ;
    11'b01000111110  : y = 8'b00111001 ;
    11'b01000111111  : y = 8'b00111001 ;
    11'b01001000000  : y = 8'b00111001 ;
    11'b01001000001  : y = 8'b00111001 ;
    11'b01001000010  : y = 8'b00111001 ;
    11'b01001000011  : y = 8'b00111001 ;
    11'b01001000100  : y = 8'b00111001 ;
    11'b01001000101  : y = 8'b00111001 ;
    11'b01001000110  : y = 8'b00111001 ;
    11'b01001000111  : y = 8'b00111001 ;
    11'b01001001000  : y = 8'b00111001 ;
    11'b01001001001  : y = 8'b00111001 ;
    11'b01001001010  : y = 8'b00111001 ;
    11'b01001001011  : y = 8'b00111001 ;
    11'b01001001100  : y = 8'b00111001 ;
    11'b01001001101  : y = 8'b00111001 ;
    11'b01001001110  : y = 8'b00111001 ;
    11'b01001001111  : y = 8'b00111001 ;
    11'b01001010000  : y = 8'b00111001 ;
    11'b01001010001  : y = 8'b00111001 ;
    11'b01001010010  : y = 8'b00111001 ;
    11'b01001010011  : y = 8'b00111001 ;
    11'b01001010100  : y = 8'b00111001 ;
    11'b01001010101  : y = 8'b00111001 ;
    11'b01001010110  : y = 8'b00111001 ;
    11'b01001010111  : y = 8'b00111001 ;
    11'b01001011000  : y = 8'b00111001 ;
    11'b01001011001  : y = 8'b00111010 ;
    11'b01001011010  : y = 8'b00111010 ;
    11'b01001011011  : y = 8'b00111010 ;
    11'b01001011100  : y = 8'b00111010 ;
    11'b01001011101  : y = 8'b00111010 ;
    11'b01001011110  : y = 8'b00111010 ;
    11'b01001011111  : y = 8'b00111010 ;
    11'b01001100000  : y = 8'b00111010 ;
    11'b01001100001  : y = 8'b00111010 ;
    11'b01001100010  : y = 8'b00111010 ;
    11'b01001100011  : y = 8'b00111010 ;
    11'b01001100100  : y = 8'b00111010 ;
    11'b01001100101  : y = 8'b00111010 ;
    11'b01001100110  : y = 8'b00111010 ;
    11'b01001100111  : y = 8'b00111010 ;
    11'b01001101000  : y = 8'b00111010 ;
    11'b01001101001  : y = 8'b00111010 ;
    11'b01001101010  : y = 8'b00111010 ;
    11'b01001101011  : y = 8'b00111010 ;
    11'b01001101100  : y = 8'b00111010 ;
    11'b01001101101  : y = 8'b00111010 ;
    11'b01001101110  : y = 8'b00111010 ;
    11'b01001101111  : y = 8'b00111010 ;
    11'b01001110000  : y = 8'b00111010 ;
    11'b01001110001  : y = 8'b00111010 ;
    11'b01001110010  : y = 8'b00111010 ;
    11'b01001110011  : y = 8'b00111010 ;
    11'b01001110100  : y = 8'b00111010 ;
    11'b01001110101  : y = 8'b00111010 ;
    11'b01001110110  : y = 8'b00111010 ;
    11'b01001110111  : y = 8'b00111010 ;
    11'b01001111000  : y = 8'b00111010 ;
    11'b01001111001  : y = 8'b00111010 ;
    11'b01001111010  : y = 8'b00111010 ;
    11'b01001111011  : y = 8'b00111010 ;
    11'b01001111100  : y = 8'b00111010 ;
    11'b01001111101  : y = 8'b00111010 ;
    11'b01001111110  : y = 8'b00111010 ;
    11'b01001111111  : y = 8'b00111010 ;
    11'b01010000000  : y = 8'b00111011 ;
    11'b01010000001  : y = 8'b00111011 ;
    11'b01010000010  : y = 8'b00111011 ;
    11'b01010000011  : y = 8'b00111011 ;
    11'b01010000100  : y = 8'b00111011 ;
    11'b01010000101  : y = 8'b00111011 ;
    11'b01010000110  : y = 8'b00111011 ;
    11'b01010000111  : y = 8'b00111011 ;
    11'b01010001000  : y = 8'b00111011 ;
    11'b01010001001  : y = 8'b00111011 ;
    11'b01010001010  : y = 8'b00111011 ;
    11'b01010001011  : y = 8'b00111011 ;
    11'b01010001100  : y = 8'b00111011 ;
    11'b01010001101  : y = 8'b00111011 ;
    11'b01010001110  : y = 8'b00111011 ;
    11'b01010001111  : y = 8'b00111011 ;
    11'b01010010000  : y = 8'b00111011 ;
    11'b01010010001  : y = 8'b00111011 ;
    11'b01010010010  : y = 8'b00111011 ;
    11'b01010010011  : y = 8'b00111011 ;
    11'b01010010100  : y = 8'b00111011 ;
    11'b01010010101  : y = 8'b00111011 ;
    11'b01010010110  : y = 8'b00111011 ;
    11'b01010010111  : y = 8'b00111011 ;
    11'b01010011000  : y = 8'b00111011 ;
    11'b01010011001  : y = 8'b00111011 ;
    11'b01010011010  : y = 8'b00111011 ;
    11'b01010011011  : y = 8'b00111011 ;
    11'b01010011100  : y = 8'b00111011 ;
    11'b01010011101  : y = 8'b00111011 ;
    11'b01010011110  : y = 8'b00111011 ;
    11'b01010011111  : y = 8'b00111011 ;
    11'b01010100000  : y = 8'b00111011 ;
    11'b01010100001  : y = 8'b00111011 ;
    11'b01010100010  : y = 8'b00111011 ;
    11'b01010100011  : y = 8'b00111011 ;
    11'b01010100100  : y = 8'b00111011 ;
    11'b01010100101  : y = 8'b00111011 ;
    11'b01010100110  : y = 8'b00111011 ;
    11'b01010100111  : y = 8'b00111011 ;
    11'b01010101000  : y = 8'b00111011 ;
    11'b01010101001  : y = 8'b00111100 ;
    11'b01010101010  : y = 8'b00111100 ;
    11'b01010101011  : y = 8'b00111100 ;
    11'b01010101100  : y = 8'b00111100 ;
    11'b01010101101  : y = 8'b00111100 ;
    11'b01010101110  : y = 8'b00111100 ;
    11'b01010101111  : y = 8'b00111100 ;
    11'b01010110000  : y = 8'b00111100 ;
    11'b01010110001  : y = 8'b00111100 ;
    11'b01010110010  : y = 8'b00111100 ;
    11'b01010110011  : y = 8'b00111100 ;
    11'b01010110100  : y = 8'b00111100 ;
    11'b01010110101  : y = 8'b00111100 ;
    11'b01010110110  : y = 8'b00111100 ;
    11'b01010110111  : y = 8'b00111100 ;
    11'b01010111000  : y = 8'b00111100 ;
    11'b01010111001  : y = 8'b00111100 ;
    11'b01010111010  : y = 8'b00111100 ;
    11'b01010111011  : y = 8'b00111100 ;
    11'b01010111100  : y = 8'b00111100 ;
    11'b01010111101  : y = 8'b00111100 ;
    11'b01010111110  : y = 8'b00111100 ;
    11'b01010111111  : y = 8'b00111100 ;
    11'b01011000000  : y = 8'b00111100 ;
    11'b01011000001  : y = 8'b00111100 ;
    11'b01011000010  : y = 8'b00111100 ;
    11'b01011000011  : y = 8'b00111100 ;
    11'b01011000100  : y = 8'b00111100 ;
    11'b01011000101  : y = 8'b00111100 ;
    11'b01011000110  : y = 8'b00111100 ;
    11'b01011000111  : y = 8'b00111100 ;
    11'b01011001000  : y = 8'b00111100 ;
    11'b01011001001  : y = 8'b00111100 ;
    11'b01011001010  : y = 8'b00111100 ;
    11'b01011001011  : y = 8'b00111100 ;
    11'b01011001100  : y = 8'b00111100 ;
    11'b01011001101  : y = 8'b00111100 ;
    11'b01011001110  : y = 8'b00111100 ;
    11'b01011001111  : y = 8'b00111100 ;
    11'b01011010000  : y = 8'b00111100 ;
    11'b01011010001  : y = 8'b00111100 ;
    11'b01011010010  : y = 8'b00111100 ;
    11'b01011010011  : y = 8'b00111100 ;
    11'b01011010100  : y = 8'b00111100 ;
    11'b01011010101  : y = 8'b00111101 ;
    11'b01011010110  : y = 8'b00111101 ;
    11'b01011010111  : y = 8'b00111101 ;
    11'b01011011000  : y = 8'b00111101 ;
    11'b01011011001  : y = 8'b00111101 ;
    11'b01011011010  : y = 8'b00111101 ;
    11'b01011011011  : y = 8'b00111101 ;
    11'b01011011100  : y = 8'b00111101 ;
    11'b01011011101  : y = 8'b00111101 ;
    11'b01011011110  : y = 8'b00111101 ;
    11'b01011011111  : y = 8'b00111101 ;
    11'b01011100000  : y = 8'b00111101 ;
    11'b01011100001  : y = 8'b00111101 ;
    11'b01011100010  : y = 8'b00111101 ;
    11'b01011100011  : y = 8'b00111101 ;
    11'b01011100100  : y = 8'b00111101 ;
    11'b01011100101  : y = 8'b00111101 ;
    11'b01011100110  : y = 8'b00111101 ;
    11'b01011100111  : y = 8'b00111101 ;
    11'b01011101000  : y = 8'b00111101 ;
    11'b01011101001  : y = 8'b00111101 ;
    11'b01011101010  : y = 8'b00111101 ;
    11'b01011101011  : y = 8'b00111101 ;
    11'b01011101100  : y = 8'b00111101 ;
    11'b01011101101  : y = 8'b00111101 ;
    11'b01011101110  : y = 8'b00111101 ;
    11'b01011101111  : y = 8'b00111101 ;
    11'b01011110000  : y = 8'b00111101 ;
    11'b01011110001  : y = 8'b00111101 ;
    11'b01011110010  : y = 8'b00111101 ;
    11'b01011110011  : y = 8'b00111101 ;
    11'b01011110100  : y = 8'b00111101 ;
    11'b01011110101  : y = 8'b00111101 ;
    11'b01011110110  : y = 8'b00111101 ;
    11'b01011110111  : y = 8'b00111101 ;
    11'b01011111000  : y = 8'b00111101 ;
    11'b01011111001  : y = 8'b00111101 ;
    11'b01011111010  : y = 8'b00111101 ;
    11'b01011111011  : y = 8'b00111101 ;
    11'b01011111100  : y = 8'b00111101 ;
    11'b01011111101  : y = 8'b00111101 ;
    11'b01011111110  : y = 8'b00111101 ;
    11'b01011111111  : y = 8'b00111101 ;
    11'b01100000000  : y = 8'b00111101 ;
    11'b01100000001  : y = 8'b00111101 ;
    11'b01100000010  : y = 8'b00111101 ;
    11'b01100000011  : y = 8'b00111101 ;
    11'b01100000100  : y = 8'b00111110 ;
    11'b01100000101  : y = 8'b00111110 ;
    11'b01100000110  : y = 8'b00111110 ;
    11'b01100000111  : y = 8'b00111110 ;
    11'b01100001000  : y = 8'b00111110 ;
    11'b01100001001  : y = 8'b00111110 ;
    11'b01100001010  : y = 8'b00111110 ;
    11'b01100001011  : y = 8'b00111110 ;
    11'b01100001100  : y = 8'b00111110 ;
    11'b01100001101  : y = 8'b00111110 ;
    11'b01100001110  : y = 8'b00111110 ;
    11'b01100001111  : y = 8'b00111110 ;
    11'b01100010000  : y = 8'b00111110 ;
    11'b01100010001  : y = 8'b00111110 ;
    11'b01100010010  : y = 8'b00111110 ;
    11'b01100010011  : y = 8'b00111110 ;
    11'b01100010100  : y = 8'b00111110 ;
    11'b01100010101  : y = 8'b00111110 ;
    11'b01100010110  : y = 8'b00111110 ;
    11'b01100010111  : y = 8'b00111110 ;
    11'b01100011000  : y = 8'b00111110 ;
    11'b01100011001  : y = 8'b00111110 ;
    11'b01100011010  : y = 8'b00111110 ;
    11'b01100011011  : y = 8'b00111110 ;
    11'b01100011100  : y = 8'b00111110 ;
    11'b01100011101  : y = 8'b00111110 ;
    11'b01100011110  : y = 8'b00111110 ;
    11'b01100011111  : y = 8'b00111110 ;
    11'b01100100000  : y = 8'b00111110 ;
    11'b01100100001  : y = 8'b00111110 ;
    11'b01100100010  : y = 8'b00111110 ;
    11'b01100100011  : y = 8'b00111110 ;
    11'b01100100100  : y = 8'b00111110 ;
    11'b01100100101  : y = 8'b00111110 ;
    11'b01100100110  : y = 8'b00111110 ;
    11'b01100100111  : y = 8'b00111110 ;
    11'b01100101000  : y = 8'b00111110 ;
    11'b01100101001  : y = 8'b00111110 ;
    11'b01100101010  : y = 8'b00111110 ;
    11'b01100101011  : y = 8'b00111110 ;
    11'b01100101100  : y = 8'b00111110 ;
    11'b01100101101  : y = 8'b00111110 ;
    11'b01100101110  : y = 8'b00111110 ;
    11'b01100101111  : y = 8'b00111110 ;
    11'b01100110000  : y = 8'b00111110 ;
    11'b01100110001  : y = 8'b00111110 ;
    11'b01100110010  : y = 8'b00111110 ;
    11'b01100110011  : y = 8'b00111110 ;
    11'b01100110100  : y = 8'b00111110 ;
    11'b01100110101  : y = 8'b00111111 ;
    11'b01100110110  : y = 8'b00111111 ;
    11'b01100110111  : y = 8'b00111111 ;
    11'b01100111000  : y = 8'b00111111 ;
    11'b01100111001  : y = 8'b00111111 ;
    11'b01100111010  : y = 8'b00111111 ;
    11'b01100111011  : y = 8'b00111111 ;
    11'b01100111100  : y = 8'b00111111 ;
    11'b01100111101  : y = 8'b00111111 ;
    11'b01100111110  : y = 8'b00111111 ;
    11'b01100111111  : y = 8'b00111111 ;
    11'b01101000000  : y = 8'b00111111 ;
    11'b01101000001  : y = 8'b00111111 ;
    11'b01101000010  : y = 8'b00111111 ;
    11'b01101000011  : y = 8'b00111111 ;
    11'b01101000100  : y = 8'b00111111 ;
    11'b01101000101  : y = 8'b00111111 ;
    11'b01101000110  : y = 8'b00111111 ;
    11'b01101000111  : y = 8'b00111111 ;
    11'b01101001000  : y = 8'b00111111 ;
    11'b01101001001  : y = 8'b00111111 ;
    11'b01101001010  : y = 8'b00111111 ;
    11'b01101001011  : y = 8'b00111111 ;
    11'b01101001100  : y = 8'b00111111 ;
    11'b01101001101  : y = 8'b00111111 ;
    11'b01101001110  : y = 8'b00111111 ;
    11'b01101001111  : y = 8'b00111111 ;
    11'b01101010000  : y = 8'b00111111 ;
    11'b01101010001  : y = 8'b00111111 ;
    11'b01101010010  : y = 8'b00111111 ;
    11'b01101010011  : y = 8'b00111111 ;
    11'b01101010100  : y = 8'b00111111 ;
    11'b01101010101  : y = 8'b00111111 ;
    11'b01101010110  : y = 8'b00111111 ;
    11'b01101010111  : y = 8'b00111111 ;
    11'b01101011000  : y = 8'b00111111 ;
    11'b01101011001  : y = 8'b00111111 ;
    11'b01101011010  : y = 8'b00111111 ;
    11'b01101011011  : y = 8'b00111111 ;
    11'b01101011100  : y = 8'b00111111 ;
    11'b01101011101  : y = 8'b00111111 ;
    11'b01101011110  : y = 8'b00111111 ;
    11'b01101011111  : y = 8'b00111111 ;
    11'b01101100000  : y = 8'b00111111 ;
    11'b01101100001  : y = 8'b00111111 ;
    11'b01101100010  : y = 8'b00111111 ;
    11'b01101100011  : y = 8'b00111111 ;
    11'b01101100100  : y = 8'b00111111 ;
    11'b01101100101  : y = 8'b00111111 ;
    11'b01101100110  : y = 8'b00111111 ;
    11'b01101100111  : y = 8'b00111111 ;
    11'b01101101000  : y = 8'b00111111 ;
    11'b01101101001  : y = 8'b00111111 ;
    11'b01101101010  : y = 8'b00111111 ;
    11'b01101101011  : y = 8'b00111111 ;
    11'b01101101100  : y = 8'b00111111 ;
    11'b01101101101  : y = 8'b00111111 ;
    11'b01101101110  : y = 8'b00111111 ;
    11'b01101101111  : y = 8'b00111111 ;
    11'b01101110000  : y = 8'b00111111 ;
    11'b01101110001  : y = 8'b00111111 ;
    11'b01101110010  : y = 8'b00111111 ;
    11'b01101110011  : y = 8'b00111111 ;
    11'b01101110100  : y = 8'b00111111 ;
    11'b01101110101  : y = 8'b00111111 ;
    11'b01101110110  : y = 8'b00111111 ;
    11'b01101110111  : y = 8'b00111111 ;
    11'b01101111000  : y = 8'b00111111 ;
    11'b01101111001  : y = 8'b00111111 ;
    11'b01101111010  : y = 8'b00111111 ;
    11'b01101111011  : y = 8'b00111111 ;
    11'b01101111100  : y = 8'b00111111 ;
    11'b01101111101  : y = 8'b00111111 ;
    11'b01101111110  : y = 8'b00111111 ;
    11'b01101111111  : y = 8'b00111111 ;
    11'b01110000000  : y = 8'b00111111 ;
    11'b01110000001  : y = 8'b00111111 ;
    11'b01110000010  : y = 8'b00111111 ;
    11'b01110000011  : y = 8'b00111111 ;
    11'b01110000100  : y = 8'b00111111 ;
    11'b01110000101  : y = 8'b00111111 ;
    11'b01110000110  : y = 8'b00111111 ;
    11'b01110000111  : y = 8'b00111111 ;
    11'b01110001000  : y = 8'b00111111 ;
    11'b01110001001  : y = 8'b00111111 ;
    11'b01110001010  : y = 8'b00111111 ;
    11'b01110001011  : y = 8'b00111111 ;
    11'b01110001100  : y = 8'b00111111 ;
    11'b01110001101  : y = 8'b00111111 ;
    11'b01110001110  : y = 8'b00111111 ;
    11'b01110001111  : y = 8'b00111111 ;
    11'b01110010000  : y = 8'b00111111 ;
    11'b01110010001  : y = 8'b00111111 ;
    11'b01110010010  : y = 8'b00111111 ;
    11'b01110010011  : y = 8'b00111111 ;
    11'b01110010100  : y = 8'b00111111 ;
    11'b01110010101  : y = 8'b00111111 ;
    11'b01110010110  : y = 8'b00111111 ;
    11'b01110010111  : y = 8'b00111111 ;
    11'b01110011000  : y = 8'b00111111 ;
    11'b01110011001  : y = 8'b00111111 ;
    11'b01110011010  : y = 8'b00111111 ;
    11'b01110011011  : y = 8'b00111111 ;
    11'b01110011100  : y = 8'b00111111 ;
    11'b01110011101  : y = 8'b00111111 ;
    11'b01110011110  : y = 8'b00111111 ;
    11'b01110011111  : y = 8'b00111111 ;
    11'b01110100000  : y = 8'b00111111 ;
    11'b01110100001  : y = 8'b00111111 ;
    11'b01110100010  : y = 8'b00111111 ;
    11'b01110100011  : y = 8'b00111111 ;
    11'b01110100100  : y = 8'b00111111 ;
    11'b01110100101  : y = 8'b00111111 ;
    11'b01110100110  : y = 8'b00111111 ;
    11'b01110100111  : y = 8'b00111111 ;
    11'b01110101000  : y = 8'b00111111 ;
    11'b01110101001  : y = 8'b00111111 ;
    11'b01110101010  : y = 8'b00111111 ;
    11'b01110101011  : y = 8'b00111111 ;
    11'b01110101100  : y = 8'b00111111 ;
    11'b01110101101  : y = 8'b00111111 ;
    11'b01110101110  : y = 8'b00111111 ;
    11'b01110101111  : y = 8'b00111111 ;
    11'b01110110000  : y = 8'b00111111 ;
    11'b01110110001  : y = 8'b00111111 ;
    11'b01110110010  : y = 8'b00111111 ;
    11'b01110110011  : y = 8'b00111111 ;
    11'b01110110100  : y = 8'b00111111 ;
    11'b01110110101  : y = 8'b00111111 ;
    11'b01110110110  : y = 8'b00111111 ;
    11'b01110110111  : y = 8'b00111111 ;
    11'b01110111000  : y = 8'b00111111 ;
    11'b01110111001  : y = 8'b00111111 ;
    11'b01110111010  : y = 8'b00111111 ;
    11'b01110111011  : y = 8'b00111111 ;
    11'b01110111100  : y = 8'b00111111 ;
    11'b01110111101  : y = 8'b00111111 ;
    11'b01110111110  : y = 8'b00111111 ;
    11'b01110111111  : y = 8'b00111111 ;
    11'b01111000000  : y = 8'b00111111 ;
    11'b01111000001  : y = 8'b00111111 ;
    11'b01111000010  : y = 8'b00111111 ;
    11'b01111000011  : y = 8'b00111111 ;
    11'b01111000100  : y = 8'b00111111 ;
    11'b01111000101  : y = 8'b00111111 ;
    11'b01111000110  : y = 8'b00111111 ;
    11'b01111000111  : y = 8'b00111111 ;
    11'b01111001000  : y = 8'b00111111 ;
    11'b01111001001  : y = 8'b00111111 ;
    11'b01111001010  : y = 8'b00111111 ;
    11'b01111001011  : y = 8'b00111111 ;
    11'b01111001100  : y = 8'b00111111 ;
    11'b01111001101  : y = 8'b00111111 ;
    11'b01111001110  : y = 8'b00111111 ;
    11'b01111001111  : y = 8'b00111111 ;
    11'b01111010000  : y = 8'b00111111 ;
    11'b01111010001  : y = 8'b00111111 ;
    11'b01111010010  : y = 8'b00111111 ;
    11'b01111010011  : y = 8'b00111111 ;
    11'b01111010100  : y = 8'b00111111 ;
    11'b01111010101  : y = 8'b00111111 ;
    11'b01111010110  : y = 8'b00111111 ;
    11'b01111010111  : y = 8'b00111111 ;
    11'b01111011000  : y = 8'b00111111 ;
    11'b01111011001  : y = 8'b00111111 ;
    11'b01111011010  : y = 8'b00111111 ;
    11'b01111011011  : y = 8'b00111111 ;
    11'b01111011100  : y = 8'b00111111 ;
    11'b01111011101  : y = 8'b00111111 ;
    11'b01111011110  : y = 8'b00111111 ;
    11'b01111011111  : y = 8'b00111111 ;
    11'b01111100000  : y = 8'b00111111 ;
    11'b01111100001  : y = 8'b00111111 ;
    11'b01111100010  : y = 8'b00111111 ;
    11'b01111100011  : y = 8'b00111111 ;
    11'b01111100100  : y = 8'b00111111 ;
    11'b01111100101  : y = 8'b00111111 ;
    11'b01111100110  : y = 8'b00111111 ;
    11'b01111100111  : y = 8'b00111111 ;
    11'b01111101000  : y = 8'b00111111 ;
    11'b01111101001  : y = 8'b00111111 ;
    11'b01111101010  : y = 8'b00111111 ;
    11'b01111101011  : y = 8'b00111111 ;
    11'b01111101100  : y = 8'b00111111 ;
    11'b01111101101  : y = 8'b00111111 ;
    11'b01111101110  : y = 8'b00111111 ;
    11'b01111101111  : y = 8'b00111111 ;
    11'b01111110000  : y = 8'b00111111 ;
    11'b01111110001  : y = 8'b00111111 ;
    11'b01111110010  : y = 8'b00111111 ;
    11'b01111110011  : y = 8'b00111111 ;
    11'b01111110100  : y = 8'b00111111 ;
    11'b01111110101  : y = 8'b00111111 ;
    11'b01111110110  : y = 8'b00111111 ;
    11'b01111110111  : y = 8'b00111111 ;
    11'b01111111000  : y = 8'b00111111 ;
    11'b01111111001  : y = 8'b00111111 ;
    11'b01111111010  : y = 8'b00111111 ;
    11'b01111111011  : y = 8'b00111111 ;
    11'b01111111100  : y = 8'b00111111 ;
    11'b01111111101  : y = 8'b00111111 ;
    11'b01111111110  : y = 8'b00111111 ;
    11'b01111111111  : y = 8'b00111111 ;
	default : y = 8'b11111111;
	endcase
end
endmodule